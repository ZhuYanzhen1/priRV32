module priRV32_IFU( 
    input clk_in,
    input rst_n,
    input [31:0] imm_decoded,
    input [4:0] rs1_decoded,
    input [4:0] rs2_decoded,
    input [4:0] rd_decoded
);



endmodule
