module decoder(
	input clk,
	input rst_n,
	output pc_address
);

endmodule
