module decoder(
	input clk,
	input rst_n,
	output [31:0] pc_address,
	input [31:0] source_data
);

endmodule
